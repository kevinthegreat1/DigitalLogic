library verilog;
use verilog.vl_types.all;
entity BinaryCounter_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        T               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end BinaryCounter_vlg_sample_tst;
