library verilog;
use verilog.vl_types.all;
entity DLatchWaveform_vlg_vec_tst is
end DLatchWaveform_vlg_vec_tst;
