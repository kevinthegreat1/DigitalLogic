library verilog;
use verilog.vl_types.all;
entity TFlipFlop_vlg_vec_tst is
end TFlipFlop_vlg_vec_tst;
