library verilog;
use verilog.vl_types.all;
entity DFlipFlop_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        D               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end DFlipFlop_vlg_sample_tst;
