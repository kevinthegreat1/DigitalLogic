module DLatchWaveform(input D, input E, output Q, output Qbar);
	DLatchKevin(D, E, Q, Qbar);
endmodule