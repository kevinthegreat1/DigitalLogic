library verilog;
use verilog.vl_types.all;
entity Thunderbird_vlg_vec_tst is
end Thunderbird_vlg_vec_tst;
