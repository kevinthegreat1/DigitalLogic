library verilog;
use verilog.vl_types.all;
entity SRNorLatch_vlg_vec_tst is
end SRNorLatch_vlg_vec_tst;
