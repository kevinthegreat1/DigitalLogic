library verilog;
use verilog.vl_types.all;
entity BasicBehavioralVerilog_vlg_vec_tst is
end BasicBehavioralVerilog_vlg_vec_tst;
