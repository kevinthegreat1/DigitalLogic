library verilog;
use verilog.vl_types.all;
entity BinaryCounter_vlg_vec_tst is
end BinaryCounter_vlg_vec_tst;
