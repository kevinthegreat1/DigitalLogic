library verilog;
use verilog.vl_types.all;
entity DFlipFlop_vlg_vec_tst is
end DFlipFlop_vlg_vec_tst;
