library verilog;
use verilog.vl_types.all;
entity ThunderbirdTest_vlg_vec_tst is
end ThunderbirdTest_vlg_vec_tst;
