library verilog;
use verilog.vl_types.all;
entity Elevator_vlg_vec_tst is
end Elevator_vlg_vec_tst;
